`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:16:41 06/18/2021 
// Design Name: 
// Module Name:    mux 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
  module mux
  #(parameter N = 32)
  (
   input wire [N-1:0] a, b,
	input wire s,
	output wire [N-1:0] out      
	);
   assign out = (s)? b : a;

  endmodule
